// You can insert code here by setting file_header_inc in file common.tpl

//=============================================================================
// Project  : generated_tb
//
// File Name: IF_sequencer.sv
//
//
// Version:   1.0
//
// Code created by Easier UVM Code Generator version 2016-08-11 on Mon Nov  5 13:07:21 2018
//=============================================================================
// Description: Sequencer for IF
//=============================================================================

`ifndef IF_SEQUENCER_SV
`define IF_SEQUENCER_SV

// Sequencer class is specialization of uvm_sequencer
typedef uvm_sequencer #(if_trans) IF_sequencer_t;


`endif // IF_SEQUENCER_SV

