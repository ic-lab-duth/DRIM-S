//register status defines
`define IDLE 2'b00
`define LANE_OPERATION 2'b01
`define STORE 2'b10
`define LOAD 2'b11

//mem state defines
`define MEM_AVAILABLE 2'b00
`define MEM_STORE 2'b01
`define MEM_LOAD 2'b10

//alu state defines
`define ALU_AVAILABLE 1'b0
`define ALU_UNAVAILABLE 1'b1
